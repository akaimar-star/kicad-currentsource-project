.title KiCad schematic
.include "../../libs/spice/THAT320-quad.lib"
.include "../../libs/spice/1N4446.lib"
.include "../../libs/spice/2N7000.REV0.lib"
.include "../../libs/spice/FQD17P06.lib"
.include "../../libs/spice/LMx58_LM2904.lib"

.param TEMP=27

*C4 GND Net-_C4-Pad2_ CAP
*C3 GND Net-_C3-Pad2_ CAP
*C1 Net-_C1-Pad1_ GND CAP
*C2 Net-_C2-Pad1_ GND CAP
XU1 Net-_U1-Pad1_ Net-_Q3-Pad3_ +15V_1 Net-_C1-Pad1_ +15V_1 Net-_Q3-Pad3_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad8_ +15V_1 Net-_C3-Pad2_ +15V_1 Net-_Q3-Pad3_ Net-_U1-Pad14_ THAT320
XU2 Net-_Q3-Pad1_ Net-_R1-Pad1_ Net-_U1-Pad1_ Net-_C2-Pad1_ Net-_U1-Pad7_ Net-_R1-Pad1_ Net-_D1-PadA_ Net-_R1-Pad1_ Net-_R1-Pad1_ Net-_U1-Pad8_ Net-_C4-Pad2_ Net-_U1-Pad14_ Net-_R1-Pad1_ Net-_D2-PadA_ THAT320
Rsafety1 Net-_D1-PadC_ GND 1k
Rload1 Net-_D2-PadC_ GND 1k
R1 Net-_R1-Pad1_ GND 20k
R2 Net-_Q3-Pad4_ GND 20k
Rset1 Net-_Q4-Pad3_ GND 330
XQ4 Net-_Q3-Pad1_ Net-_Q4-Pad2_ Net-_Q4-Pad3_ 2N7000
XU3 Net-_U3-Pad3_ Net-_Q4-Pad3_ +15V_1 GND Net-_Q4-Pad2_ LM358
Vref1 Net-_U3-Pad3_ GND 3.3
Vsource1 +15V_1 GND 15
XQ3 Net-_Q3-Pad4_ Net-_Q3-Pad1_ Net-_Q3-Pad3_ FQD17P06
D1 Net-_D1-PadA_ Net-_D1-PadC_ 1N4446
D2 Net-_D2-PadA_ Net-_D2-PadC_ 1N4446


.options savecurrents
.save @Rload1[i]
.save @Rsafety1[i]


* Control Statements 
.control
run
parameter sweep
* resistive divider, R1 swept from start_r to stop_r
let start_r = 0
let stop_r = 3k
let delta_r = 100
let r_act = start_r
let iload=unitvec(stop_r/delta_r+1)
let Rload=unitvec(stop_r/delta_r+1)
let isafety=unitvec(stop_r/delta_r+1)
let iideal=unitvec(stop_r/delta_r+1)
* loop
while r_act le stop_r
  alter Rload1 r_act
  op
  let iload[r_act/delta_r]=$&@Rload1[i]
  let isafety[r_act/delta_r]=$&@Rsafety1[i]
  let iideal[r_act/delta_r]=10m
  let Rload[r_act/delta_r]=$&r_act
  let r_act = r_act + delta_r
end

settype current iload
settype current isafety
settype current iideal
settype res-sweep Rload
plot iload isafety iideal vs 'Rload'
.endc
.end
